`define initial_read 3'd0
`define M0_AR_S0 3'd1
`define M0_AR_S1 3'd2
`define M0_read 3'd3
`define M1_AR_S1 3'd4
`define M1_AR_S0 3'd5
`define M1_read 3'd6


`define initial_write 3'd0
`define M1_AW_S1 3'd1
`define M1_write_S1 3'd2
`define M1_AW_S0 3'd3
`define M1_write_S0 3'd4
`define M1_RESP 3'd5

