`define initial_read 4'd0
`define M0_AR_S0 4'd1
`define M0_AR_S1 4'd2
`define M0_AR_S2 4'd3
`define M0_AR_S4 4'd4
`define M0_read 4'd5
`define M1_AR_S0 4'd6
`define M1_AR_S1 4'd7
`define M1_AR_S2 4'd8
`define M1_AR_S4 4'd9
`define M1_read 4'd10



`define initial_write 3'd0
`define M1_write_S1 3'd1
`define M1_write_S2 3'd2
`define M1_write_S4 3'd3
`define M1_RESP 3'd4

